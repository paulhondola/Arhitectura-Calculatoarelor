module ex2(

);


endmodule